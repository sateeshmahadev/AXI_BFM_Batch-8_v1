`ifndef FIFO_BFM_32B_WR_INCR_ALLIGNED_TEST_AWLEN_12_TO_15_INCLUDED_
`define FIFO_BFM_32B_WR_INCR_ALLIGNED_TEST_AWLEN_12_TO_15_INCLUDED_

//-----------------------------------------------------------------------------
// Class: fifo_bfm_32b_wr_incr_alligned_test_awlen_12_to_15 
// Description of the class:
// This class provides the test case for fifo_bfm_32b_wr_incr_alligned_awlen_12_to_15 
// where awlenn can be in the range [12, 15]
//-----------------------------------------------------------------------------
class fifo_bfm_32b_wr_incr_alligned_test_awlen_12_to_15 extends fifo_base_test;
  `uvm_component_utils(fifo_bfm_32b_wr_incr_alligned_test_awlen_12_to_15)

  //Local variables of this test through which we send values to the sequence
  bit[31:0] wdata_seq[$];
  bit[3:0] awlenn;
  bit[31:0] addr;
  bit[3:0] wstrbb = 4'hf;
  bit[1:0] awburstt = 1;
  bit[2:0] awsizee = 2;

  // Sequence handles for write transactions
  fifo_bfm_wr_incr_alligned_sequence fifo_bfm_wr_incr_alligned_sequence_h;  //write fifo sequence
  axi4_slave_nbk_write_32b_transfer_seq axi4_slave_nbk_write_32b_transfer_seq_h; //wr response sequence by avip slave

  //-----------------------------------------------------------------------------
  // Constructor: new
  // Initializes the fifo_bfm_32b_wr_incr_alligned_test_awlen_12_to_15 class object
  //
  // Parameters:
  //  name - instance name of the fifo_bfm_32b_wr_incr_alligned_test_awlen_12_to_15 
  //  parent - parent under which this component is created
  //-----------------------------------------------------------------------------
  function new(string name = "fifo_bfm_32b_wr_incr_alligned_test_awlen_12_to_15", uvm_component parent = null);
    super.new(name, parent);
    // Randomize awlenn within the range [12, 15]
    void'(std::randomize(awlenn) with {awlenn inside {[12:15]};});
    `uvm_info("UVM_TEST", $sformatf("AWLEN = %h", awlenn), UVM_MEDIUM)
    void'(std::randomize(addr) with {addr % ((2**awsizee) * 8) == 0;});
    `uvm_info("UVM_TEST", $sformatf("Address = %h", addr), UVM_MEDIUM)
    void'(std::randomize(wdata_seq) with {wdata_seq.size() == awlenn + 1;});
  endfunction

  //-----------------------------------------------------------------------------
  // Function: build_phase
  // Creates the required sequences
  //
  // Parameters:
  //  phase - stores the current phase 
  //-----------------------------------------------------------------------------
  function void build_phase(uvm_phase phase);
    super.build_phase(phase);
    axi4_slave_nbk_write_32b_transfer_seq_h = axi4_slave_nbk_write_32b_transfer_seq::type_id::create("axi4_slave_nbk_write_32b_transfer_seq_h");
    fifo_bfm_wr_incr_alligned_sequence_h = fifo_bfm_wr_incr_alligned_sequence::type_id::create("fifo_bfm_wr_incr_alligned_sequence_h");
  endfunction

  //-----------------------------------------------------------------------------
  // Task: run_phase
  // Assign values from local variables of test to the sequence variables and starts the two sequences
  //
  // Parameters:
  //  phase - stores the current phase 
  //-----------------------------------------------------------------------------
  task run_phase(uvm_phase phase);
    `uvm_info(get_type_name(), $sformatf("fifo_bfm_32b_wr_incr_alligned_test_awlen_12_to_15"), UVM_LOW)

    phase.raise_objection(this);

    // Configure the write sequence parameters through local variables of test
    fifo_bfm_wr_incr_alligned_sequence_h.awlenn = awlenn;
    fifo_bfm_wr_incr_alligned_sequence_h.addr = addr;
    fifo_bfm_wr_incr_alligned_sequence_h.wstrbb = wstrbb;
    fifo_bfm_wr_incr_alligned_sequence_h.awburstt = awburstt;
    fifo_bfm_wr_incr_alligned_sequence_h.awsizee = awsizee;
    fifo_bfm_wr_incr_alligned_sequence_h.wdata_seq = wdata_seq;
   
    // Start the write sequence and the avip write response sequence concurrently
    fork
      begin
        forever begin
          axi4_slave_nbk_write_32b_transfer_seq_h.start(env_h.axi_slave_agent_h.axi4_slave_write_seqr_h);
        end
      end
    join_none

    // Start the FIFO write sequence
    fifo_bfm_wr_incr_alligned_sequence_h.start(env_h.write_fifo_agent_h.write_fifo_sequencer_h);

    phase.drop_objection(this);
  endtask
endclass
`endif

